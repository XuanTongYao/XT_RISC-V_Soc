//----------内存RAM----------//
`define INST_RAM_DEPTH 512
`define INST_RAM_ADDR_WIDTH $clog2(`INST_RAM_DEPTH * 4)
`define RAM_DEPTH 512
`define RAM_ADDR_WIDTH $clog2(`RAM_DEPTH * 4)

`define INST_RAM_LEN (`INST_RAM_DEPTH*4)
`define DATA_RAM_LEN (`RAM_DEPTH*4)
`define INST_RAM_BASE 0
`define DATA_RAM_BASE (`INST_RAM_BASE+`INST_RAM_LEN)


//----------XT_HB总线----------//

// 外设占用地址长度
`define DOMAIN_XT_HB_LEN 32
`define DOMAIN_WISHBONE_LEN 256
`define DOMAIN_XT_LB_LEN 256

// 外设地址偏移定义
`define DOMAIN_XT_HB_OFFSET 0
`define DOMAIN_WISHBONE_OFFSET (`DOMAIN_XT_HB_OFFSET+`DOMAIN_XT_HB_LEN)
`define DOMAIN_XT_LB_OFFSET (`DOMAIN_WISHBONE_OFFSET+`DOMAIN_WISHBONE_LEN)

// 外设基地址定义
`define BUS_DOMAIN_BASE (`DATA_RAM_BASE+`DATA_RAM_LEN)
`define DOMAIN_XT_HB_BASE (`BUS_DOMAIN_BASE+`DOMAIN_XT_HB_OFFSET)
`define DOMAIN_WISHBONE_BASE (`BUS_DOMAIN_BASE+`DOMAIN_WISHBONE_OFFSET)
`define DOMAIN_XT_LB_BASE (`BUS_DOMAIN_BASE+`DOMAIN_XT_LB_OFFSET)
