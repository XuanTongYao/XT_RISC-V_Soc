
//----------XT_HB总线----------//

// 外设占用地址长度
`define DEBUG_LEN 4
`define EINT_CTRL_LEN 8
`define SYSTEM_TIMER_LEN 16
`define UART_LEN 4
`define WISHBONE_LEN 256
`define XT_LB_LEN 256

// 外设地址偏移定义
`define DEBUG_OFFSET 0
`define EINT_CTRL_OFFSET (`DEBUG_OFFSET+`DEBUG_LEN)
`define SYSTEM_TIMER_OFFSET (`EINT_CTRL_OFFSET+`EINT_CTRL_LEN)
`define UART_OFFSET (`SYSTEM_TIMER_OFFSET+`SYSTEM_TIMER_LEN)
`define WISHBONE_OFFSET (`UART_OFFSET+`UART_LEN)
`define XT_LB_OFFSET (`WISHBONE_OFFSET+`WISHBONE_LEN)

// 外设基地址定义
`define PERIPHERALS_BASE (`DATA_RAM_BASE+`DATA_RAM_LEN)
`define DEBUG_BASE (`PERIPHERALS_BASE+`DEBUG_OFFSET)
`define EINT_CTRL_BASE (`PERIPHERALS_BASE+`EINT_CTRL_OFFSET)
`define SYSTEM_TIMER_BASE (`PERIPHERALS_BASE+`SYSTEM_TIMER_OFFSET)
`define UART_BASE (`PERIPHERALS_BASE+`UART_OFFSET)
`define WISHBONE_BASE (`PERIPHERALS_BASE+`WISHBONE_OFFSET)
`define XT_LB_BASE (`PERIPHERALS_BASE+`XT_LB_OFFSET)


//----------WISHBONE总线----------//
// 外设占用地址长度
`define FLASH_LEN 5

// 外设地址偏移定义
`define FLASH_OFFSET 32'h70

// 外设基地址定义
`define FLASH_BASE (`WISHBONE_BASE+`FLASH_OFFSET)

