package Utils_Pkg;


  // 读写片选
  typedef struct packed {
    logic ren;
    logic wen;
  } sel_t;



endpackage
