// 0:使能寄存器  4:待处理中断寄存器
module External_INT_Ctrl
  import Utils_Pkg::sel_t;
  import SystemPeripheral_Pkg::*;
#(
    parameter int INT_NUM = 32
) (
    input rst_sync,
    input hb_clk,
    input sys_peripheral_t sys_share,
    input sel_t sel,
    output logic [31:0] rdata,

    input [INT_NUM-1:0] irq_source,
    // 自定义中断代码，用于向量跳转，大于等于16的部分，只有27位，原来的代码最长也只有31位
    output logic [26:0] custom_int_code,
    output logic mextern_int

);

  logic [INT_NUM-1:0] INT_enable_reg;
  logic [INT_NUM-1:0] INT_pending_reg;
  always_ff @(posedge hb_clk) begin
    if (rst_sync) begin
      INT_enable_reg  <= 0;
      INT_pending_reg <= 0;
    end else begin
      if (sel.wen && sys_share.waddr == 'd0) begin
        INT_enable_reg <= sys_share.wdata[INT_NUM-1:0];
      end
      INT_pending_reg <= irq_source & INT_enable_reg;
    end
  end


  logic [5:0] int_id;
  always_comb begin
    int id;
    id = 0;
    int_id = 0;
    for (int i = 0; i < INT_NUM; ++i) begin
      if (INT_pending_reg[i]) begin
        id = i + 1;
        int_id = id[5:0];
        break;
      end
    end
    mextern_int = |INT_pending_reg;
    custom_int_code = {21'b0, int_id};
  end



  // 总线读
  always_ff @(posedge hb_clk) begin
    if (sel.ren) begin
      if (sys_share.raddr == 'd0) begin
        rdata <= INT_enable_reg;
      end else begin
        rdata <= INT_pending_reg;
      end
    end
  end


endmodule
