//----------异常原因代码定义----------//


`define EXCEPTION_INVALID_INST 4'd2
`define EXCEPTION_EBREAK 4'd3
`define EXCEPTION_MECALL 4'd11

